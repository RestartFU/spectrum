module internal

pub const ascii = "HxNjF7upSSAFZkDENZKduZ8JhXBXmLwmL7pPxYY6B8UzQMAPMUZt6Xa4XDETzx9UpCCUGQ1xs18oNse2XzB8faeP4opZ4NCp6Ur4j7w4BHcLuspBAGvPh5mA5Hyhd5Ppdy4XLfFF75ffvUciaHjRiCC9QeMsfuXwouZshSRZiQgferDRqUi6XpvG82WEr4UjATtDkkRK16eFhVcX3WCpkp23cDLGKLyitqU7hut3MHhmv2o2vwnxm7uN4UYqXoAYK3VYkd"
