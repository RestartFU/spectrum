module command

pub interface Valuable {
	value() string
}