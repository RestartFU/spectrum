module packet

pub enum ID {
	handshake
	login
	hwid_check
	hwid_check_result
	message_data
}
